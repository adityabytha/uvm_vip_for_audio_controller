




class i2s_sequencer extends uvm_sequencer#(i2s_tx);
	`uvm_component_utils(i2s_sequencer)
	`NEW
endclass
