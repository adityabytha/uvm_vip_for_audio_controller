




class dac_sequencer extends uvm_sequencer#(dac_tx);
	`uvm_component_utils(dac_sequencer)
	`NEW
endclass
