




class spdif_sequencer extends uvm_sequencer#(spdif_tx);
	`uvm_component_utils(spdif_sequencer)
	`NEW
endclass
