




class main_sequencer extends uvm_sequencer#(audio_tx);
	`uvm_component_utils(main_sequencer)
	`NEW
endclass
